library verilog;
use verilog.vl_types.all;
entity TestB_Control is
end TestB_Control;
