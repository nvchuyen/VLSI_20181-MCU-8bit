library verilog;
use verilog.vl_types.all;
entity TestB_Instruction is
end TestB_Instruction;
