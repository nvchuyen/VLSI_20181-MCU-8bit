library verilog;
use verilog.vl_types.all;
entity TestB_Register is
end TestB_Register;
