library verilog;
use verilog.vl_types.all;
entity TestB_PC is
end TestB_PC;
