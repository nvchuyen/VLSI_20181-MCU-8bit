library verilog;
use verilog.vl_types.all;
entity TestB_InPutOP is
end TestB_InPutOP;
