library verilog;
use verilog.vl_types.all;
entity TestB_MCU is
end TestB_MCU;
